-- Copyright (C) 2017  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 17.1.0 Build 590 10/25/2017 SJ Lite Edition"
-- CREATED		"Tue Mar 03 10:06:27 2020"

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.ALL;  

-- Add the library and use clauses before the design unit declaration
library altera; 
use altera.altera_primitives_components.all;

LIBRARY work;


ENTITY ROM_READER_V2 IS 
	PORT
	(
		TRIGGER_IN :  IN  STD_LOGIC;
		CLK :  IN  STD_LOGIC;
		RESET :  IN  STD_LOGIC;
		READ_ENA :  OUT  STD_LOGIC;
		ROM_ADDR :  OUT  STD_LOGIC_VECTOR(9 DOWNTO 0);
		SOP	: OUT STD_LOGIC; --FIRST SAMPLE OUT
		EOP	:	OUT STD_LOGIC --SECONDS SAMPLE OUT
	);
END ROM_READER_V2;

ARCHITECTURE rtl OF ROM_READER_V2 IS 

SIGNAL	RESETn :  STD_LOGIC;
SIGNAL	SOP_OUT : STD_LOGIC;	--WIRES
SIGNAL 	EOP_OUT	: STD_LOGIC; --WIRES
SIGNAL	Q_OUT : STD_LOGIC_VECTOR(9 DOWNTO 0);
SIGNAL	COUNTER : NATURAL;
signal	read_ena_out : std_logic;
signal	dff1:	std_logic;
signal	dff0: std_logic;
signal	cnt_ena_ff: std_logic;
signal	cout : std_logic;

	


BEGIN 
	
		--COUNTER <=  to_integer(unsigned(Q_OUT));
		--my_slv <= std_logic_vector(to_unsigned(my_int, my_slv'length));
		
		Q_OUT <= std_logic_vector(to_unsigned(COUNTER, 10));
		
		SOP <= SOP_OUT;
		EOP <= EOP_OUT;
		
		READ_ENA <= cnt_ena_ff;
		ROM_ADDR <= Q_OUT;

		
	
		
	--10bitcounter
	process (CLK,RESET,cnt_ena_ff)
		variable cnt : natural range 0 to 1023 := 0;
	begin
				
		if (rising_edge(clk)) then
		
				if (RESET = '1') then
				-- Reset the counter to 0
				cnt := 0;

				elsif cnt_ena_ff = '1' then		
				
					--reset counter
					if cnt = 1023 then
					cnt := 0;
					else
					-- Increment the counter if counting is enabled			   
					cnt := cnt + 1;
					end if;
					
				
				end if;
				
		end if;

		-- Output the current count
		COUNTER <= cnt;
		
		-- some AND gates
		if ( cnt = 0 and cnt_ena_ff = '1') then
			SOP_OUT <= '1';
		else
			SOP_OUT <= '0';
		end if;
		
		if (cnt = 1023 and cnt_ena_ff = '1') then
			EOP_OUT <= '1';
			cout <= '1';
		else
			EOP_OUT <= '0';
			cout <= '0';
		end if;
		
		--Q_OUT <= std_logic_vector(to_unsigned(cnt, 10));
	end process;

	

--TRIGGER_IN CAPTURE
--dff0	
	process(RESET, TRIGGER_IN, dff1)
begin
	if((RESET = '1') or (dff1 = '1')) then
		dff0 <= '0';
	elsif (rising_edge(TRIGGER_IN)) then
		dff0 <= '1';
	end if;
end process;

--dff1
process (CLK)
begin
	if (rising_edge(CLK)) then
		dff1 <= dff0;
	end if;
end process;

--cnt_ena_ff
process(CLK, dff1, cout, reset)
begin
	if(reset = '1') then
		cnt_ena_ff <= '0';
	elsif ((dff1 = '1') or (cout = '1')) then
		if (rising_edge(CLK)) then
			cnt_ena_ff <= dff1;
		end if;
	end if;
end process;

	
	
RESETn <= NOT(RESET);	

END rtl;